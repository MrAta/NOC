`ifndef _noc_params_vh_
`define _noc_params_vh_

	`define conn_entries 16
	`define num_credit_delay 5
	`define num_of_vcs 6
	`define max_cycles 100000
	`define num_of_routers 4
	`define vcs_size 3

`endif
